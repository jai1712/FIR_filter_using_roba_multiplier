module adder(a,b,sum);
input [63:0]a,b;
output [63:0]sum;

assign sum=a+b;

endmodule